module Hexadecimalto7Seg(A, D);

input [3:0] A;
output reg [6:0] D;

always @(A)
begin
    case (A)
        0: D[6:0] = 7'b1000000;  // 0
        1: D[6:0]  = 7'b1111001;  // 1
        2: D[6:0]  = 7'b0100100;  // 2
        3: D[6:0]  = 7'b0110000;  // 3
        4: D[6:0]  = 7'b0011001;  // 4
        5: D[6:0]  = 7'b0010010;  // 5
        6: D[6:0]  = 7'b0000010;  // 6
        7: D[6:0]  = 7'b1111000;  // 7
        8: D[6:0]  = 7'b0000000;  // 8
        9: D[6:0]  = 7'b0010000;
		  10: D[6:0]  = 7'b0001000;
		  11: D[6:0]  = 7'b0000011;
		  12: D[6:0]  = 7'b1000110;
		  13: D[6:0]  = 7'b0100001;	
		  14: D[6:0]  = 7'b0000110;
		  15: D[6:0]  = 7'b0001110;			
        default: D[6:0]  = 7'b0111111;  // Default (blank or error)
    endcase
end



endmodule

